
module on_chip_memory #(
	parameter IP_TYPE 		= "OCM",
	parameter IP_VERSION 	= 32'h1, 
	parameter IP_ID 		= 32'h4c60de2
)
(
    input  wire    [9:0] addr_A,
    input  wire   [17:0] din_A,
    input  wire    [9:0] addr_B,
    input  wire          wen_A,
    input  wire          ren_B,
    output wire   [17:0] dout_B,
    input  wire          clk
);


//------------------------------------------------------------------------------
// Signals
//------------------------------------------------------------------------------

wire          sys_clk;
wire    [9:0] addr_A_1;
wire    [9:0] addr_B_1;
wire   [17:0] din_A_1;
wire   [17:0] dout_B_1;
wire          wen_A_1;
wire          ren_B_1;
wire   [15:0] bram_out_B;
wire    [1:0] rparity_B;

//------------------------------------------------------------------------------
// Combinatorial Logic
//------------------------------------------------------------------------------

assign addr_A_1 = addr_A;
assign din_A_1 = din_A;
assign addr_B_1 = addr_B;
assign wen_A_1 = wen_A;
assign ren_B_1 = ren_B;
assign dout_B = dout_B_1;
assign sys_clk = clk;
assign dout_B_1[17:0] = {rparity_B[1], bram_out_B[15:8], rparity_B[0], bram_out_B[7:0]};

TDP_RAM18KX2 # (
    .INIT1({16384{1'b0}}),
    .INIT1_PARITY({2048{1'b0}}),
    .WRITE_WIDTH_A1(18),
    .READ_WIDTH_B1(18)
  )
  TDP_RAM18KX2_inst (
    .WEN_A1(wen_A_1),
    .REN_B1(ren_B_1),
    .CLK_A1(clk),
    .CLK_B1(clk),
    .BE_A1({2{1'd1}}),
    .ADDR_A1({addr_A_1[9:0], {4{1'd0}}}),
    .ADDR_B1({addr_B_1[9:0], {4{1'd0}}}),
    .WDATA_A1({din_A_1[16:9], din_A_1[7:0]}),
    .WPARITY_A1({din_A_1[17], din_A_1[8]}),
    .RDATA_B1(bram_out_B[15:0]),
    .RPARITY_B1(rparity_B[1:0])
  );

endmodule

// -----------------------------------------------------------------------------
//  Auto-Generated by LiteX on 2024-06-12 12:51:12.
//------------------------------------------------------------------------------

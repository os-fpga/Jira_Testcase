`define Total_instances 1
module ram_inst_sp_36 #(parameter AWIDTH = 10, DWIDTH = 36) (
  input clock0, we,
  input [AWIDTH-1:0] addr, 
  input [DWIDTH-1:0] din,
  input [$clog2(`Total_instances)-1:0] id, 
  output [DWIDTH-1:0] dout);

parameter [80:0] MODE_BITS =81'h0;

wire [DWIDTH-1:0] dout_arr [0:`Total_instances-1];
reg [`Total_instances-1:0] we_arr;
wire [DWIDTH-1:0] open_wire1 [0:`Total_instances-1];
genvar i;

generate
  for (i=0;i<`Total_instances;i=i+1) begin
    RS_TDP36K  #(.MODE_BITS(MODE_BITS))
      inst1(
    .ADDR_A1({ addr, 5'h00 }),
    .ADDR_A2({ addr[8:0], 5'h00 }),
    .ADDR_B1(0),
    .ADDR_B2(0),
    .BE_A1(3),
    .BE_A2(3),
    .BE_B1(3),
    .BE_B2(3),
    .CLK_A1(clock0),
    .CLK_A2(clock0),
    .CLK_B1(clock0),
    .CLK_B2(clock0),
    .FLUSH1(0),
    .FLUSH2(0),
    .RDATA_A1({dout_arr[i][33:32],dout_arr[i][15:0]}),
    .RDATA_A2({dout_arr[i][35:34],dout_arr[i][31:16]}),
    .RDATA_B1(),
    .RDATA_B2(),
    .REN_A1(~we_arr[i]),
    .REN_A2(~we_arr[i]),
    .REN_B1(0),
    .REN_B2(0),
    .WDATA_A1({din[33:32],din[15:0]}),
    .WDATA_A2({din[35:34],din[31:16]}),
    .WDATA_B1(0),
    .WDATA_B2(0),
    .WEN_A1(we_arr[i]),
    .WEN_A2(we_arr[i]),
    .WEN_B1(0),
    .WEN_B2(0)
  );
 
end
endgenerate
 
assign dout = dout_arr[id];

integer j;

always @ (*) begin
  for(j=0;j<`Total_instances;j=j+1)begin
    we_arr[j] = 'd0;
  end
    we_arr[id] = we;
end

endmodule

/* Generated by Yosys 0.18+10 (git sha1 2b3815b19, gcc 9.4.0 -fPIC -Os) */

// (* top =  1  *)
// (* src = "/nfs_scratch/scratch/CompilerValidation/abdul_hameed/reggression/Compiler_Validation/RTL_testcases/Memory_Designs/Simple_dual_port_rams/ram_simple_dp_dc_512x32/rtl/ram_simple_dp_dc_512x32.v:1" *)
// module rams_sp_rwe(we, read_clock, write_clock, read_addr, write_addr, dout, din);
//   (* unused_bits = "32 33 34 35" *)
//   wire [35:0] \$auto$memory_bram.cc:844:replace_memory$48 ;
//   (* src = "/nfs_cadtools/raptor/instl_dir/bin/../share/yosys/rapidsilicon/genesis/brams_map.v:318.14-318.19" *)
//   (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35" *)
//   wire [35:0] \$techmap64\ram.0.0.0.DOBDO ;
//   (* src = "/nfs_scratch/scratch/CompilerValidation/abdul_hameed/reggression/Compiler_Validation/RTL_testcases/Memory_Designs/Simple_dual_port_rams/ram_simple_dp_dc_512x32/rtl/ram_simple_dp_dc_512x32.v:2" *)
//   input [31:0] din;
//   wire [31:0] din;
//   (* src = "/nfs_scratch/scratch/CompilerValidation/abdul_hameed/reggression/Compiler_Validation/RTL_testcases/Memory_Designs/Simple_dual_port_rams/ram_simple_dp_dc_512x32/rtl/ram_simple_dp_dc_512x32.v:5" *)
//   output [31:0] dout;
//   wire [31:0] dout;
//   (* src = "/nfs_scratch/scratch/CompilerValidation/abdul_hameed/reggression/Compiler_Validation/RTL_testcases/Memory_Designs/Simple_dual_port_rams/ram_simple_dp_dc_512x32/rtl/ram_simple_dp_dc_512x32.v:3" *)
//   input [8:0] read_addr;
//   wire [8:0] read_addr;
//   (* src = "/nfs_scratch/scratch/CompilerValidation/abdul_hameed/reggression/Compiler_Validation/RTL_testcases/Memory_Designs/Simple_dual_port_rams/ram_simple_dp_dc_512x32/rtl/ram_simple_dp_dc_512x32.v:4" *)
//   input read_clock;
//   wire read_clock;
//   (* src = "/nfs_scratch/scratch/CompilerValidation/abdul_hameed/reggression/Compiler_Validation/RTL_testcases/Memory_Designs/Simple_dual_port_rams/ram_simple_dp_dc_512x32/rtl/ram_simple_dp_dc_512x32.v:4" *)
//   input we;
//   wire we;
//   (* src = "/nfs_scratch/scratch/CompilerValidation/abdul_hameed/reggression/Compiler_Validation/RTL_testcases/Memory_Designs/Simple_dual_port_rams/ram_simple_dp_dc_512x32/rtl/ram_simple_dp_dc_512x32.v:3" *)
//   input [8:0] write_addr;
//   wire [8:0] write_addr;
//   (* src = "/nfs_scratch/scratch/CompilerValidation/abdul_hameed/reggression/Compiler_Validation/RTL_testcases/Memory_Designs/Simple_dual_port_rams/ram_simple_dp_dc_512x32/rtl/ram_simple_dp_dc_512x32.v:4" *)
//   input write_clock;
//   wire write_clock;
//   (* module_not_derived = 32'h00000001 *)
//   (* src = "/nfs_cadtools/raptor/instl_dir/bin/../share/yosys/rapidsilicon/genesis/brams_map.v:408.9-442.3" *)
//   RS_TDP36K #(
//     .MODE_BITS(81'h00140281b6c0140140db6)
//   ) \ram.0.0.0  (
//     .ADDR_A1({ 1'h0, read_addr, 5'h00 }),
//     .ADDR_A2({ read_addr, 5'h00 }),
//     .ADDR_B1({ 1'h0, write_addr, 5'h00 }),
//     .ADDR_B2({ write_addr, 5'h00 }),
//     .BE_A1(2'h3),
//     .BE_A2(2'h3),
//     .BE_B1({ we, we }),
//     .BE_B2({ we, we }),
//     .CLK_A1(read_clock),
//     .CLK_A2(read_clock),
//     .CLK_B1(write_clock),
//     .CLK_B2(write_clock),
//     .FLUSH1(1'h0),
//     .FLUSH2(1'h0),
//     .RDATA_A1(dout[17:0]),
//     .RDATA_A2({ \$auto$memory_bram.cc:844:replace_memory$48 [35:32], dout[31:18] }),
//     .RDATA_B1(\$techmap64\ram.0.0.0.DOBDO [17:0]),
//     .RDATA_B2(\$techmap64\ram.0.0.0.DOBDO [35:18]),
//     .REN_A1(1'h1),
//     .REN_A2(1'h1),
//     .REN_B1(1'h0),
//     .REN_B2(1'h0),
//     .WDATA_A1(18'h3ffff),
//     .WDATA_A2(18'h3ffff),
//     .WDATA_B1(din[17:0]),
//     .WDATA_B2({ 4'hx, din[31:18] }),
//     .WEN_A1(1'h0),
//     .WEN_A2(1'h0),
//     .WEN_B1(we),
//     .WEN_B2(we)
//   );
//   assign \$auto$memory_bram.cc:844:replace_memory$48 [31:0] = dout;
// endmodule

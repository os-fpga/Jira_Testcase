module test(a,b);

    input wire a;
    output reg b;

    assign b = a;

endmodule